name=Namn
email=Email
mobileNr=Mobilnr
password=Lösenord
location=Plats
date=Datum
information=Information
creator=Skapare